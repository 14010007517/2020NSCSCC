`timescale 1 ns / 1 ps

module cpu_core (
    
);
    

    
endmodule